`define DATA_WIDTH 5
