// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

module debug_array();

    logic [3:0] test_a;

    logic test_b [3:0];

endmodule
