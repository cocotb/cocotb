module debug_array;

    // Equivalent to std_logic_vector(3 downto 0)
    logic [3:0] test_a;

    // Equivalent to array (3 downto 0) of std_logic
    logic test_b [3:0];

endmodule
