-- Copyright cocotb contributors
-- Licensed under the Revised BSD License, see LICENSE for details.
-- SPDX-License-Identifier: BSD-3-Clause

use work.cocotb_package_pkg_1.all;
use work.cocotb_package_pkg_2.all;

entity cocotb_package is
end entity cocotb_package;

architecture test of cocotb_package is
    constant seven_int : integer := 7;
begin
end architecture test;
