-- Copyright cocotb contributors
-- Licensed under the Revised BSD License, see LICENSE for details.
-- SPDX-License-Identifier: BSD-3-Clause

package integers_pkg is
    subtype my_integer is integer range -100 to 100;
end package integers_pkg;
