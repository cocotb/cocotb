module issue_3239
    (input union packed {
           logic [3:0] a;
           logic [1:0][1:0] b;
     } t);
endmodule : issue_3239
