// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

`timescale 1us/1us

module test (
    input logic KPFIVTM1LHY0OFUNXF0XZO1RV535NNU4A8QWR12BLQXJ98PMM1P552QC0T089PUJPB4POUJZLBS19S8XNMPGJV2QK3AJUW98X7RU56ZV4IMFIPDJI81E5B9HNW94Q9APLMMK3VPHS1VB1QVPQDG7VOTLY2NT3F4080OUXSC68H0JZF7KQ0O6GGN3DARXC03CSZL7TE6B7R47366SB54T5Q4MOR5BT3L5S0S3NM8MALXPHZKCUA6AR5U391GGDYG5LB7JGKAHSIREODSNGW7FAYNRTTXFFCRL4U3ZQA6DH1RKCFKGDG9WMF81IX5YSAINQSP14F2FJV0GYEM3R4LUFFSWOZKK5MGKS25RLROJFEQDC8L2XY07728MM7V516ZXH1YFS0AL1GPLH03N5EL0RQVY61EVEQEJCYDT0ZBBN1ZLC5BDQU83NF8N953MU6A99SDNPCTSOD2W9WY69ZL64JHURFHA5DT7KQC7T4KASR5CAG85ONU3F2XWYA97JHDN9V9SBS39MYMYERJ338O6JQYCHX7SH8FB2VL2PI7DOQWB3NXTA8CQM7YKT34L6U3O42WWMI7NHKUIBO4U9MBP176000FU39WET32RG4PHLYYGWFMKPYPCUFE46RFSQDELLXU31ZZH0OJCGEFUDR2USDUYZ3XPBQ6RC0XARPG2Z1GHCESILHJOF7503PHKWUKDVM2V18WB16CB7AAQ8C4C6E7FXUB3E89Q0ZJSKQFYNZPSKYKGXURV3V5C0SHU9QQ2GFUTP38ORCSWN0QYIX9H0SKJEXPC5U1D3QN9PRT0QPOVM7H5EGQ4E449YTSHUMJW1TT2S6EVIPPIR9ZMFCOWPYXRSNJEQ3OCKGDUW2ZX2AS7N5GBUY7NOAR2P7BK5YPOA6APVAH12V86V2YQZ2M56HLNAD785GI4GMFSCI5P3LNFM0CLSBUEJXCVT695N5D3GC8T0HKAN0BZDV1ZMI0WZ3QUVABNYFOJHXXBUW5OK5MQ46NMK3W0FMCKWVPP6265,
    output logic o);

assign o = KPFIVTM1LHY0OFUNXF0XZO1RV535NNU4A8QWR12BLQXJ98PMM1P552QC0T089PUJPB4POUJZLBS19S8XNMPGJV2QK3AJUW98X7RU56ZV4IMFIPDJI81E5B9HNW94Q9APLMMK3VPHS1VB1QVPQDG7VOTLY2NT3F4080OUXSC68H0JZF7KQ0O6GGN3DARXC03CSZL7TE6B7R47366SB54T5Q4MOR5BT3L5S0S3NM8MALXPHZKCUA6AR5U391GGDYG5LB7JGKAHSIREODSNGW7FAYNRTTXFFCRL4U3ZQA6DH1RKCFKGDG9WMF81IX5YSAINQSP14F2FJV0GYEM3R4LUFFSWOZKK5MGKS25RLROJFEQDC8L2XY07728MM7V516ZXH1YFS0AL1GPLH03N5EL0RQVY61EVEQEJCYDT0ZBBN1ZLC5BDQU83NF8N953MU6A99SDNPCTSOD2W9WY69ZL64JHURFHA5DT7KQC7T4KASR5CAG85ONU3F2XWYA97JHDN9V9SBS39MYMYERJ338O6JQYCHX7SH8FB2VL2PI7DOQWB3NXTA8CQM7YKT34L6U3O42WWMI7NHKUIBO4U9MBP176000FU39WET32RG4PHLYYGWFMKPYPCUFE46RFSQDELLXU31ZZH0OJCGEFUDR2USDUYZ3XPBQ6RC0XARPG2Z1GHCESILHJOF7503PHKWUKDVM2V18WB16CB7AAQ8C4C6E7FXUB3E89Q0ZJSKQFYNZPSKYKGXURV3V5C0SHU9QQ2GFUTP38ORCSWN0QYIX9H0SKJEXPC5U1D3QN9PRT0QPOVM7H5EGQ4E449YTSHUMJW1TT2S6EVIPPIR9ZMFCOWPYXRSNJEQ3OCKGDUW2ZX2AS7N5GBUY7NOAR2P7BK5YPOA6APVAH12V86V2YQZ2M56HLNAD785GI4GMFSCI5P3LNFM0CLSBUEJXCVT695N5D3GC8T0HKAN0BZDV1ZMI0WZ3QUVABNYFOJHXXBUW5OK5MQ46NMK3W0FMCKWVPP6265;

endmodule
