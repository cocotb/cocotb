parameter DATA_BYTES = 8;