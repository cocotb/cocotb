`define DATA_LAST 64
