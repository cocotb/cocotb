// This file is public domain, it can be freely copied without restrictions.
// SPDX-License-Identifier: CC0-1.0

import cds_rnm_pkg::*;

package nettypes_pkg;

  nettype wreal1driver voltage_net;

endpackage
