// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

`timescale 1 ps / 1 ps

module top (
    input logic placeholder
);

endmodule
