// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause


module cocotb_initial;

    int foo;
    initial foo = 123;

endmodule
