// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

/* verilator public_on */
package cocotb_package_pkg_1;
    parameter int five_int = 5;
    parameter logic [31:0] eight_logic = 8;
    parameter logic [63:0] long_param = '1;
endpackage

package cocotb_package_pkg_2;
    parameter int eleven_int = 11;
endpackage

parameter int unit_four_int = 4;

/* verilator public_off */
