`define DATA_LAST 3
