`define DATA_BYTES 8
