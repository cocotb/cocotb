package cocotb_package_pkg_1;
    parameter int five_int = 5;
    parameter logic [31:0] eight_logic = 8;
endpackage

package cocotb_package_pkg_2;
    parameter int eleven_int = 11;
endpackage

parameter int unit_four_int = 4;
