// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

module debug_array;

    reg [3:0] test_a;

    initial begin
        test_a   = 4'b0000;
    end

endmodule
