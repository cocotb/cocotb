-- This file is public domain, it can be freely copied without restrictions.
-- SPDX-License-Identifier: CC0-1.0

entity dummy is
end dummy;

architecture empty of dummy is
begin
end empty;
