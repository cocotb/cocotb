// Copyright cocotb contributors
// Licensed under the Revised BSD License, see LICENSE for details.
// SPDX-License-Identifier: BSD-3-Clause

`timescale 1us/1us

interface sv_if();
  logic a;
  reg b;
  wire c;
endinterface

module top ();

sv_if sv_if_i();

sv_if sv_if_arr[3]();

endmodule
