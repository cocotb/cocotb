parameter DATA_LAST = 64;