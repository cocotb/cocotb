parameter DATA_WIDTH = 32;