module debug_array;

    logic [3:0] test_a;

    logic test_b [3:0];

endmodule
